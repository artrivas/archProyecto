module mainfsm (
	clk,
	reset,
	Op,
	Funct,
	Branch,
	MemtoReg,
	MemW,
	ALUSrc,
	ImmSrc,
	RegW,
	RegSrc,
	Branch,
	ALUOp
);
	input wire clk;
	input wire reset;
	input wire [1:0] Op;
	input wire [5:0] Funct;
	output wire Branch;
	output wire MemtoReg;
	output wire MemW;
	output wire ALUSrc;
	output wire [1:0] ImmSrc;
	output wire RegW;
	output wire [1:0] RegSrc;
	output wire Branch;
	output wire ALUOp;
	reg [3:0] state;
	reg [3:0] nextstate;
	reg [12:0] controls;

	localparam [3:0] FETCH = 0;
	localparam [3:0] DECODE = 1;
	localparam [3:0] MEMADR = 2;
	localparam [3:0] MEMREAD = 3;
	localparam [3:0] MEMWB = 4;
	localparam [3:0] MEMWRITE = 5;
	localparam [3:0] EXECUTER = 6;
	localparam [3:0] EXECUTEI = 7;
	localparam [3:0] ALUWB = 8;
	localparam [3:0] BRANCH = 9;
	localparam [3:0] UNKNOWN = 10;

	// state register
	always @(posedge clk or posedge reset)
		if (reset)
			state <= FETCH;
		else
			state <= nextstate;
	

	// ADD CODE BELOW
  	// Finish entering the next state logic below.  We've completed the 
  	// first two states, FETCH and DECODE, for you.

  	// next state logic
	always @(*)
		casex (state)
			FETCH: nextstate = DECODE;
			DECODE:
				case (Op)
					2'b00:
						if (Funct[5])
							nextstate = EXECUTEI;
						else
							nextstate = EXECUTER;
					2'b01: nextstate = MEMADR;
					2'b10: nextstate = BRANCH;
					default: nextstate = UNKNOWN;
				endcase
			MEMADR: 
                case (Funct[0])
                    1'b0:
                        nextstate = MEMWRITE;
                    1'b1:
                        nextstate = MEMREAD;
                endcase
			MEMREAD: nextstate = MEMWB;
			EXECUTER: nextstate = ALUWB;
			EXECUTEI: nextstate = ALUWB;
			default: nextstate = FETCH;
		endcase

	// ADD CODE BELOW
	// Finish entering the output logic below.  We've entered the
	// output logic for the first two states, FETCH and DECODE, for you.

	// state-dependent output logic
	always @(*)
		case (state)
			FETCH: controls = 12'b000101001100;
			DECODE: controls = 12'b000001001100;
			EXECUTER: controls = 12'b000000000001;
			EXECUTEI: controls = 12'b000000000011; 
			ALUWB: controls = 12'b001000000000; 
			MEMADR: controls = 12'b000000000010; 
			MEMWRITE:controls = 12'b010010000000; 
			MEMREAD: controls = 12'b000010000000; 
			MEMWB: controls = 12'b001000100000; 
			BRANCH: controls = 12'b100001010010;
			default: controls = 12'bxxxxxxxxxxxx;
		endcase
	assign {Branch, MemtoReg, MemW, ALUSrc, ImmSrc, RegW, RegSrc, Branch, ALUSrcB, ALUOp} = controls;
endmodule